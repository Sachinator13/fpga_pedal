module counter(
	input clk,
	output [3:0] count
);


endmodule