module counter(
	input clk,
	output [15:0] count
);


endmodule